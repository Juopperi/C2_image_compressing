library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all; 
use IEEE.STD_LOGIC_TEXTIO.ALL;


entity quantization_tb is
end quantization_tb;

architecture test of quantization_tb is
  component quantization
    port (
        clk    : in std_logic;
        Y   : in  std_logic_vector (1023 downto 0); 
        Cb  : in  std_logic_vector (1023 downto 0);
        Cr  : in  std_logic_vector (1023 downto 0);
        Y_out  : out std_logic_vector (1023 downto 0);
        Cb_out : out std_logic_vector (1023 downto 0);
        Cr_out : out std_logic_vector (1023 downto 0)
    );
  end component;

        signal clk    : std_logic :='0';
        signal Y_out  : std_logic_vector (1023 downto 0); 
        signal Cb_out : std_logic_vector (1023 downto 0);
        signal Cr_out : std_logic_vector (1023 downto 0);

    -- inputs from DCT (retrieved from matlab)
    signal Y : std_logic_vector (1023 downto 0):= 
        "0000000001100010" & "0010101010101010" & "0011000000100101" & "1011001010101111" & 
        "1100010000100110" & "0001010100001111" & "0001100100111101" & "1111111101000110" & 
        "0011101010101000" & "0100000100001110" & "0101101101101101" & "0010011111100100" & 
        "1111000101010111" & "0011100001010010" & "1110000011000110" & "1110010011000110" & 
        "1111101011000011" & "0111011101001111" & "0000111011010101" & "0000101100111111" & 
        "0011110000111011" & "0000000010111010" & "1101110001110101" & "0001100111111111" & 
        "0100010100111001" & "1101001001011011" & "1101010111001010" & "0001000001000011" & 
        "0100110011111111" & "1111111101111100" & "1011000111100001" & "1100010001110010" & 
        "1111100000111000" & "1101001100001011" & "0011100011001011" & "0000000011000010" & 
        "1110000001100111" & "1101001010001111" & "0000000011010001" & "0100110110010011" & 
        "1110100001100001" & "0101101010100100" & "1101001011011010" & "0100000101010110" & 
        "1111111111011000" & "1100110001011010" & "1100100001110000" & "1101001001101110" & 
        "1000010010010010" & "1110001011100001" & "0000000010000011" & "0010110001110101" & 
        "1100111101100110" & "1100010011111110" & "1100010001111011" & "1111111101011010" & 
        "1101110001110101" & "1000101001110010" & "1101000001101100" & "1101000011111100" & 
        "0000000000001101" & "1100110000000111" & "0011010000000110" & "1100111101100111";
    signal Cb :  std_logic_vector (1023 downto 0) := 
        "1100110001010111" & "1101001001111111" & "0100010100111010" & "0010100011000110" & 
        "0000001011111011" & "1111101100001000" & "1111101001100001" & "1111111010100001" & 
        "0000011000011111" & "0000110010111001" & "0000000110100100" & "0000010100001111" & 
        "1111111000111111" & "1111101011000001" & "0000001001010111" & "0000010111010111" & 
        "0001000101010110" & "1010100111000011" & "1111111111110101" & "1111111100001010" & 
        "0000001111110101" & "0000010101101000" & "1111111011010001" & "1111111100000110" & 
        "1111011000001111" & "0001100011110111" & "0000000011101100" & "0000010000101001" & 
        "1111111001010101" & "1111110111010110" & "0000001000000101" & "0000010001001100" & 
        "0000001001001110" & "0000000000111001" & "1111111001000101" & "1111111010010101" & 
        "0000001010100000" & "0000001010000101" & "1111111011000100" & "1111111000000001" & 
        "1111111111001010" & "1111101101110101" & "0000001101100010" & "0000000100011100" & 
        "1111111011010010" & "1111111010001100" & "0000000101111000" & "0000001101001001" & 
        "1111111110101011" & "0000010111101111" & "1111111000000011" & "1111111110110101" & 
        "0000000011111110" & "0000000100001011" & "1111111010110000" & "1111111101101101" & 
        "1111111011011111" & "1111111110101100" & "0000000100000100" & "0000000001110101" & 
        "1111111010001101" & "1111111110101001" & "1111111111110001" & "0000000011101011";
    signal Cr : std_logic_vector (1023 downto 0) := 
        "0101001011111111" & "0010001100111011" & "1111111110101100" & "1111111111100000" & 
        "1111111111001110" & "1111111110101101" & "1111111111011011" & "0000000000011011" & 
        "0001100001000100" & "0001001000111111" & "1111111101101001" & "1111111110100001" & 
        "1111111111000000" & "1111111111010110" & "1111111111001100" & "1111111110111001" & 
        "0001011101001001" & "1110011000110010" & "0000001100111100" & "1111111111000001" & 
        "1111111110101100" & "1111111111101111" & "0000000000010011" & "0000000100110100" & 
        "1101001100001101" & "0000001000101110" & "0001011000101100" & "1111111111100011" & 
        "0000000000101110" & "0000000000111000" & "1111111101100111" & "1111111111001110" & 
        "0000000000010011" & "0000000100001011" & "0000000100101101" & "0000000100010100" & 
        "0000000001110110" & "0000000001001101" & "0000000001001011" & "0000000001100000" & 
        "0001001000010011" & "0000000101001010" & "1111101010100000" & "0000000100111100" & 
        "0000000111100010" & "0000000101100000" & "0000000101010000" & "0000000000000001" & 
        "1111111111010001" & "0000001100001001" & "0000000111001100" & "0000000111011100" & 
        "0000000100111010" & "0000000100110001" & "0000000001011011" & "0000000001001001" & 
        "0000000100101110" & "0000000100010001" & "0000000001101000" & "0000000001001010" & 
        "0000000001110010" & "0000000000111101" & "1111111111110101" & "0000000000100001";

    file Y_file : TEXT open write_mode is "Y.txt";
    file Cb_file : TEXT open write_mode is "Cb.txt";
    file Cr_file : TEXT open write_mode is "Cr.txt";

  begin
    uut : quantization
      port map(
        clk => clk,
        Y => Y,
        Cb => Cb,
        Cr => Cr,
        Y_out => Y_out,
        Cb_out => Cb_out,
        Cr_out => Cr_out
      );

    process
    begin
        wait for 10 ns;
        clk <= not clk;
    end process;

    process
        variable L : line;
    begin
        -- Wait for some time (optional)
        wait for 2500 ns;

        -- Write vector to the file
        write(L, Y_out); 
        writeline(Y_file, L);
        write(L, Cb_out); 
        writeline(Cb_file, L);
        write(L, Cr_out); 
        writeline(Cr_file, L);

        wait; -- stop simulation
    end process;

end test;
