wire [32*64-1:0] dct_coeffs =  {
    32'h00005A82,
    32'h00005A82,
    32'h00005A82,
    32'h00005A82,
    32'h00005A82,
    32'h00005A82,
    32'h00005A82,
    32'h00005A82,
    32'h00007D8A,
    32'h00006A6D,
    32'h0000471C,
    32'h000018F8,
    32'hFFFFE708,
    32'hFFFFB8E4,
    32'hFFFF9593,
    32'hFFFF8276,
    32'h00007641,
    32'h000030FB,
    32'hFFFFCF05,
    32'hFFFF89BF,
    32'hFFFF89BF,
    32'hFFFFCF05,
    32'h000030FB,
    32'h00007641,
    32'h00006A6D,
    32'hFFFFE708,
    32'hFFFF8276,
    32'hFFFFB8E4,
    32'h0000471C,
    32'h00007D8A,
    32'h000018F8,
    32'hFFFF9593,
    32'h00005A82,
    32'hFFFFA57E,
    32'hFFFFA57E,
    32'h00005A82,
    32'h00005A82,
    32'hFFFFA57E,
    32'hFFFFA57E,
    32'h00005A82,
    32'h0000471C,
    32'hFFFF8276,
    32'h000018F8,
    32'h00006A6D,
    32'hFFFF9593,
    32'hFFFFE708,
    32'h00007D8A,
    32'hFFFFB8E4,
    32'h000030FB,
    32'hFFFF89BF,
    32'h00007641,
    32'hFFFFCF05,
    32'hFFFFCF05,
    32'h00007641,
    32'hFFFF89BF,
    32'h000030FB,
    32'h000018F8,
    32'hFFFFB8E4,
    32'h00006A6D,
    32'hFFFF8276,
    32'h00007D8A,
    32'hFFFF9593,
    32'h0000471C,
    32'hFFFFE708
};
