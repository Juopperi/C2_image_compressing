wire [32*64-1:0] dct_coeffs =  {
    32'h00005A82,
    32'h00005A82,
    32'h00005A82,
    32'h00005A82,
    32'h00005A82,
    32'h00005A82,
    32'h00005A82,
    32'h00005A82,
    32'h00007D8A,
    32'h00006A6E,
    32'h0000471D,
    32'h000018F9,
    32'hFFFFE707,
    32'hFFFFB8E3,
    32'hFFFF9592,
    32'hFFFF8276,
    32'h00007642,
    32'h000030FC,
    32'hFFFFCF04,
    32'hFFFF89BE,
    32'hFFFF89BE,
    32'hFFFFCF04,
    32'h000030FC,
    32'h00007642,
    32'h00006A6E,
    32'hFFFFE707,
    32'hFFFF8276,
    32'hFFFFB8E3,
    32'h0000471D,
    32'h00007D8A,
    32'h000018F9,
    32'hFFFF9592,
    32'h00005A82,
    32'hFFFFA57E,
    32'hFFFFA57E,
    32'h00005A82,
    32'h00005A82,
    32'hFFFFA57E,
    32'hFFFFA57E,
    32'h00005A82,
    32'h0000471D,
    32'hFFFF8276,
    32'h000018F9,
    32'h00006A6E,
    32'hFFFF9592,
    32'hFFFFE707,
    32'h00007D8A,
    32'hFFFFB8E3,
    32'h000030FC,
    32'hFFFF89BE,
    32'h00007642,
    32'hFFFFCF04,
    32'hFFFFCF04,
    32'h00007642,
    32'hFFFF89BE,
    32'h000030FC,
    32'h000018F9,
    32'hFFFFB8E3,
    32'h00006A6E,
    32'hFFFF8276,
    32'h00007D8A,
    32'hFFFF9592,
    32'h0000471D,
    32'hFFFFE707
};
