wire [32*64-1:0] luma_qtable_inv = {
    32'h00001000,
    32'h00001746,
    32'h0000199A,
    32'h00001000,
    32'h00000AAB,
    32'h00000666,
    32'h00000505,
    32'h00000432,
    32'h00001555,
    32'h00001555,
    32'h00001249,
    32'h00000D79,
    32'h000009D9,
    32'h0000046A,
    32'h00000444,
    32'h000004A8,
    32'h00001249,
    32'h000013B1,
    32'h00001000,
    32'h00000AAB,
    32'h00000666,
    32'h0000047E,
    32'h000003B6,
    32'h00000492,
    32'h00001249,
    32'h00000F0F,
    32'h00000BA3,
    32'h000008D4,
    32'h00000505,
    32'h000002F1,
    32'h00000333,
    32'h00000421,
    32'h00000E39,
    32'h00000BA3,
    32'h000006EB,
    32'h00000492,
    32'h000003C4,
    32'h00000259,
    32'h0000027C,
    32'h00000353,
    32'h00000AAB,
    32'h00000750,
    32'h000004A8,
    32'h00000400,
    32'h00000329,
    32'h00000276,
    32'h00000244,
    32'h000002C8,
    32'h00000539,
    32'h00000400,
    32'h00000348,
    32'h000002F1,
    32'h0000027C,
    32'h0000021E,
    32'h00000222,
    32'h00000289,
    32'h0000038E,
    32'h000002C8,
    32'h000002B2,
    32'h0000029D,
    32'h00000249,
    32'h0000028F,
    32'h0000027C,
    32'h00000296
};

wire [32*64-1:0] chroma_qtable_inv = {
    32'h00000F0F,
    32'h00000E39,
    32'h00000AAB,
    32'h00000572,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000E39,
    32'h00000C31,
    32'h000009D9,
    32'h000003E1,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000AAB,
    32'h000009D9,
    32'h00000492,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000572,
    32'h000003E1,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296,
    32'h00000296
};

